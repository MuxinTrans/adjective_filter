// megafunction wizard: %PARALLEL_ADD%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: parallel_add 

// ============================================================
// File Name: pAdd_80.v
// Megafunction Name(s):
// 			parallel_add
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 17.0.0 Build 595 04/25/2017 SJ Standard Edition
// ************************************************************


//Copyright (C) 2017  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Intel and sold by Intel or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module pAdd_80 (
	data0x,
	data10x,
	data11x,
	data12x,
	data13x,
	data14x,
	data15x,
	data16x,
	data17x,
	data18x,
	data19x,
	data1x,
	data20x,
	data21x,
	data22x,
	data23x,
	data24x,
	data25x,
	data26x,
	data27x,
	data28x,
	data29x,
	data2x,
	data30x,
	data31x,
	data32x,
	data33x,
	data34x,
	data35x,
	data36x,
	data37x,
	data38x,
	data39x,
	data3x,
	data40x,
	data41x,
	data42x,
	data43x,
	data44x,
	data45x,
	data46x,
	data47x,
	data48x,
	data49x,
	data4x,
	data50x,
	data51x,
	data52x,
	data53x,
	data54x,
	data55x,
	data56x,
	data57x,
	data58x,
	data59x,
	data5x,
	data60x,
	data61x,
	data62x,
	data63x,
	data64x,
	data65x,
	data66x,
	data67x,
	data68x,
	data69x,
	data6x,
	data70x,
	data71x,
	data72x,
	data73x,
	data74x,
	data75x,
	data76x,
	data77x,
	data78x,
	data79x,
	data7x,
	data8x,
	data9x,
	result);

	input	[29:0]  data0x;
	input	[29:0]  data10x;
	input	[29:0]  data11x;
	input	[29:0]  data12x;
	input	[29:0]  data13x;
	input	[29:0]  data14x;
	input	[29:0]  data15x;
	input	[29:0]  data16x;
	input	[29:0]  data17x;
	input	[29:0]  data18x;
	input	[29:0]  data19x;
	input	[29:0]  data1x;
	input	[29:0]  data20x;
	input	[29:0]  data21x;
	input	[29:0]  data22x;
	input	[29:0]  data23x;
	input	[29:0]  data24x;
	input	[29:0]  data25x;
	input	[29:0]  data26x;
	input	[29:0]  data27x;
	input	[29:0]  data28x;
	input	[29:0]  data29x;
	input	[29:0]  data2x;
	input	[29:0]  data30x;
	input	[29:0]  data31x;
	input	[29:0]  data32x;
	input	[29:0]  data33x;
	input	[29:0]  data34x;
	input	[29:0]  data35x;
	input	[29:0]  data36x;
	input	[29:0]  data37x;
	input	[29:0]  data38x;
	input	[29:0]  data39x;
	input	[29:0]  data3x;
	input	[29:0]  data40x;
	input	[29:0]  data41x;
	input	[29:0]  data42x;
	input	[29:0]  data43x;
	input	[29:0]  data44x;
	input	[29:0]  data45x;
	input	[29:0]  data46x;
	input	[29:0]  data47x;
	input	[29:0]  data48x;
	input	[29:0]  data49x;
	input	[29:0]  data4x;
	input	[29:0]  data50x;
	input	[29:0]  data51x;
	input	[29:0]  data52x;
	input	[29:0]  data53x;
	input	[29:0]  data54x;
	input	[29:0]  data55x;
	input	[29:0]  data56x;
	input	[29:0]  data57x;
	input	[29:0]  data58x;
	input	[29:0]  data59x;
	input	[29:0]  data5x;
	input	[29:0]  data60x;
	input	[29:0]  data61x;
	input	[29:0]  data62x;
	input	[29:0]  data63x;
	input	[29:0]  data64x;
	input	[29:0]  data65x;
	input	[29:0]  data66x;
	input	[29:0]  data67x;
	input	[29:0]  data68x;
	input	[29:0]  data69x;
	input	[29:0]  data6x;
	input	[29:0]  data70x;
	input	[29:0]  data71x;
	input	[29:0]  data72x;
	input	[29:0]  data73x;
	input	[29:0]  data74x;
	input	[29:0]  data75x;
	input	[29:0]  data76x;
	input	[29:0]  data77x;
	input	[29:0]  data78x;
	input	[29:0]  data79x;
	input	[29:0]  data7x;
	input	[29:0]  data8x;
	input	[29:0]  data9x;
	output	[36:0]  result;

	wire [36:0] sub_wire81;
	wire [29:0] sub_wire80 = data79x[29:0];
	wire [29:0] sub_wire79 = data78x[29:0];
	wire [29:0] sub_wire78 = data77x[29:0];
	wire [29:0] sub_wire77 = data76x[29:0];
	wire [29:0] sub_wire76 = data75x[29:0];
	wire [29:0] sub_wire75 = data74x[29:0];
	wire [29:0] sub_wire74 = data73x[29:0];
	wire [29:0] sub_wire73 = data72x[29:0];
	wire [29:0] sub_wire72 = data71x[29:0];
	wire [29:0] sub_wire71 = data70x[29:0];
	wire [29:0] sub_wire70 = data69x[29:0];
	wire [29:0] sub_wire69 = data68x[29:0];
	wire [29:0] sub_wire68 = data67x[29:0];
	wire [29:0] sub_wire67 = data66x[29:0];
	wire [29:0] sub_wire66 = data65x[29:0];
	wire [29:0] sub_wire65 = data64x[29:0];
	wire [29:0] sub_wire64 = data63x[29:0];
	wire [29:0] sub_wire63 = data62x[29:0];
	wire [29:0] sub_wire62 = data61x[29:0];
	wire [29:0] sub_wire61 = data60x[29:0];
	wire [29:0] sub_wire60 = data59x[29:0];
	wire [29:0] sub_wire59 = data58x[29:0];
	wire [29:0] sub_wire58 = data57x[29:0];
	wire [29:0] sub_wire57 = data56x[29:0];
	wire [29:0] sub_wire56 = data55x[29:0];
	wire [29:0] sub_wire55 = data54x[29:0];
	wire [29:0] sub_wire54 = data53x[29:0];
	wire [29:0] sub_wire53 = data52x[29:0];
	wire [29:0] sub_wire52 = data51x[29:0];
	wire [29:0] sub_wire51 = data50x[29:0];
	wire [29:0] sub_wire50 = data49x[29:0];
	wire [29:0] sub_wire49 = data48x[29:0];
	wire [29:0] sub_wire48 = data47x[29:0];
	wire [29:0] sub_wire47 = data46x[29:0];
	wire [29:0] sub_wire46 = data45x[29:0];
	wire [29:0] sub_wire45 = data44x[29:0];
	wire [29:0] sub_wire44 = data43x[29:0];
	wire [29:0] sub_wire43 = data42x[29:0];
	wire [29:0] sub_wire42 = data41x[29:0];
	wire [29:0] sub_wire41 = data40x[29:0];
	wire [29:0] sub_wire40 = data39x[29:0];
	wire [29:0] sub_wire39 = data38x[29:0];
	wire [29:0] sub_wire38 = data37x[29:0];
	wire [29:0] sub_wire37 = data36x[29:0];
	wire [29:0] sub_wire36 = data35x[29:0];
	wire [29:0] sub_wire35 = data34x[29:0];
	wire [29:0] sub_wire34 = data33x[29:0];
	wire [29:0] sub_wire33 = data32x[29:0];
	wire [29:0] sub_wire32 = data31x[29:0];
	wire [29:0] sub_wire31 = data30x[29:0];
	wire [29:0] sub_wire30 = data29x[29:0];
	wire [29:0] sub_wire29 = data28x[29:0];
	wire [29:0] sub_wire28 = data27x[29:0];
	wire [29:0] sub_wire27 = data26x[29:0];
	wire [29:0] sub_wire26 = data25x[29:0];
	wire [29:0] sub_wire25 = data24x[29:0];
	wire [29:0] sub_wire24 = data23x[29:0];
	wire [29:0] sub_wire23 = data22x[29:0];
	wire [29:0] sub_wire22 = data21x[29:0];
	wire [29:0] sub_wire21 = data20x[29:0];
	wire [29:0] sub_wire20 = data19x[29:0];
	wire [29:0] sub_wire19 = data18x[29:0];
	wire [29:0] sub_wire18 = data17x[29:0];
	wire [29:0] sub_wire17 = data16x[29:0];
	wire [29:0] sub_wire16 = data15x[29:0];
	wire [29:0] sub_wire15 = data14x[29:0];
	wire [29:0] sub_wire14 = data13x[29:0];
	wire [29:0] sub_wire13 = data12x[29:0];
	wire [29:0] sub_wire12 = data11x[29:0];
	wire [29:0] sub_wire11 = data10x[29:0];
	wire [29:0] sub_wire10 = data9x[29:0];
	wire [29:0] sub_wire9 = data8x[29:0];
	wire [29:0] sub_wire8 = data7x[29:0];
	wire [29:0] sub_wire7 = data6x[29:0];
	wire [29:0] sub_wire6 = data5x[29:0];
	wire [29:0] sub_wire5 = data4x[29:0];
	wire [29:0] sub_wire4 = data3x[29:0];
	wire [29:0] sub_wire3 = data2x[29:0];
	wire [29:0] sub_wire2 = data1x[29:0];
	wire [29:0] sub_wire0 = data0x[29:0];
	wire [2399:0] sub_wire1 = {sub_wire80, sub_wire79, sub_wire78, sub_wire77, sub_wire76, sub_wire75, sub_wire74, sub_wire73, sub_wire72, sub_wire71, sub_wire70, sub_wire69, sub_wire68, sub_wire67, sub_wire66, sub_wire65, sub_wire64, sub_wire63, sub_wire62, sub_wire61, sub_wire60, sub_wire59, sub_wire58, sub_wire57, sub_wire56, sub_wire55, sub_wire54, sub_wire53, sub_wire52, sub_wire51, sub_wire50, sub_wire49, sub_wire48, sub_wire47, sub_wire46, sub_wire45, sub_wire44, sub_wire43, sub_wire42, sub_wire41, sub_wire40, sub_wire39, sub_wire38, sub_wire37, sub_wire36, sub_wire35, sub_wire34, sub_wire33, sub_wire32, sub_wire31, sub_wire30, sub_wire29, sub_wire28, sub_wire27, sub_wire26, sub_wire25, sub_wire24, sub_wire23, sub_wire22, sub_wire21, sub_wire20, sub_wire19, sub_wire18, sub_wire17, sub_wire16, sub_wire15, sub_wire14, sub_wire13, sub_wire12, sub_wire11, sub_wire10, sub_wire9, sub_wire8, sub_wire7, sub_wire6, sub_wire5, sub_wire4, sub_wire3, sub_wire2, sub_wire0};
	wire [36:0] result = sub_wire81[36:0];

	parallel_add	parallel_add_component (
				.data (sub_wire1),
				.result (sub_wire81)
				// synopsys translate_off
				,
				.aclr (),
				.clken (),
				.clock ()
				// synopsys translate_on
				);
	defparam
		parallel_add_component.msw_subtract = "NO",
		parallel_add_component.pipeline = 0,
		parallel_add_component.representation = "SIGNED",
		parallel_add_component.result_alignment = "LSB",
		parallel_add_component.shift = 0,
		parallel_add_component.size = 80,
		parallel_add_component.width = 30,
		parallel_add_component.widthr = 37;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: MSW_SUBTRACT STRING "NO"
// Retrieval info: CONSTANT: PIPELINE NUMERIC "0"
// Retrieval info: CONSTANT: REPRESENTATION STRING "SIGNED"
// Retrieval info: CONSTANT: RESULT_ALIGNMENT STRING "LSB"
// Retrieval info: CONSTANT: SHIFT NUMERIC "0"
// Retrieval info: CONSTANT: SIZE NUMERIC "80"
// Retrieval info: CONSTANT: WIDTH NUMERIC "30"
// Retrieval info: CONSTANT: WIDTHR NUMERIC "37"
// Retrieval info: USED_PORT: data0x 0 0 30 0 INPUT NODEFVAL "data0x[29..0]"
// Retrieval info: USED_PORT: data10x 0 0 30 0 INPUT NODEFVAL "data10x[29..0]"
// Retrieval info: USED_PORT: data11x 0 0 30 0 INPUT NODEFVAL "data11x[29..0]"
// Retrieval info: USED_PORT: data12x 0 0 30 0 INPUT NODEFVAL "data12x[29..0]"
// Retrieval info: USED_PORT: data13x 0 0 30 0 INPUT NODEFVAL "data13x[29..0]"
// Retrieval info: USED_PORT: data14x 0 0 30 0 INPUT NODEFVAL "data14x[29..0]"
// Retrieval info: USED_PORT: data15x 0 0 30 0 INPUT NODEFVAL "data15x[29..0]"
// Retrieval info: USED_PORT: data16x 0 0 30 0 INPUT NODEFVAL "data16x[29..0]"
// Retrieval info: USED_PORT: data17x 0 0 30 0 INPUT NODEFVAL "data17x[29..0]"
// Retrieval info: USED_PORT: data18x 0 0 30 0 INPUT NODEFVAL "data18x[29..0]"
// Retrieval info: USED_PORT: data19x 0 0 30 0 INPUT NODEFVAL "data19x[29..0]"
// Retrieval info: USED_PORT: data1x 0 0 30 0 INPUT NODEFVAL "data1x[29..0]"
// Retrieval info: USED_PORT: data20x 0 0 30 0 INPUT NODEFVAL "data20x[29..0]"
// Retrieval info: USED_PORT: data21x 0 0 30 0 INPUT NODEFVAL "data21x[29..0]"
// Retrieval info: USED_PORT: data22x 0 0 30 0 INPUT NODEFVAL "data22x[29..0]"
// Retrieval info: USED_PORT: data23x 0 0 30 0 INPUT NODEFVAL "data23x[29..0]"
// Retrieval info: USED_PORT: data24x 0 0 30 0 INPUT NODEFVAL "data24x[29..0]"
// Retrieval info: USED_PORT: data25x 0 0 30 0 INPUT NODEFVAL "data25x[29..0]"
// Retrieval info: USED_PORT: data26x 0 0 30 0 INPUT NODEFVAL "data26x[29..0]"
// Retrieval info: USED_PORT: data27x 0 0 30 0 INPUT NODEFVAL "data27x[29..0]"
// Retrieval info: USED_PORT: data28x 0 0 30 0 INPUT NODEFVAL "data28x[29..0]"
// Retrieval info: USED_PORT: data29x 0 0 30 0 INPUT NODEFVAL "data29x[29..0]"
// Retrieval info: USED_PORT: data2x 0 0 30 0 INPUT NODEFVAL "data2x[29..0]"
// Retrieval info: USED_PORT: data30x 0 0 30 0 INPUT NODEFVAL "data30x[29..0]"
// Retrieval info: USED_PORT: data31x 0 0 30 0 INPUT NODEFVAL "data31x[29..0]"
// Retrieval info: USED_PORT: data32x 0 0 30 0 INPUT NODEFVAL "data32x[29..0]"
// Retrieval info: USED_PORT: data33x 0 0 30 0 INPUT NODEFVAL "data33x[29..0]"
// Retrieval info: USED_PORT: data34x 0 0 30 0 INPUT NODEFVAL "data34x[29..0]"
// Retrieval info: USED_PORT: data35x 0 0 30 0 INPUT NODEFVAL "data35x[29..0]"
// Retrieval info: USED_PORT: data36x 0 0 30 0 INPUT NODEFVAL "data36x[29..0]"
// Retrieval info: USED_PORT: data37x 0 0 30 0 INPUT NODEFVAL "data37x[29..0]"
// Retrieval info: USED_PORT: data38x 0 0 30 0 INPUT NODEFVAL "data38x[29..0]"
// Retrieval info: USED_PORT: data39x 0 0 30 0 INPUT NODEFVAL "data39x[29..0]"
// Retrieval info: USED_PORT: data3x 0 0 30 0 INPUT NODEFVAL "data3x[29..0]"
// Retrieval info: USED_PORT: data40x 0 0 30 0 INPUT NODEFVAL "data40x[29..0]"
// Retrieval info: USED_PORT: data41x 0 0 30 0 INPUT NODEFVAL "data41x[29..0]"
// Retrieval info: USED_PORT: data42x 0 0 30 0 INPUT NODEFVAL "data42x[29..0]"
// Retrieval info: USED_PORT: data43x 0 0 30 0 INPUT NODEFVAL "data43x[29..0]"
// Retrieval info: USED_PORT: data44x 0 0 30 0 INPUT NODEFVAL "data44x[29..0]"
// Retrieval info: USED_PORT: data45x 0 0 30 0 INPUT NODEFVAL "data45x[29..0]"
// Retrieval info: USED_PORT: data46x 0 0 30 0 INPUT NODEFVAL "data46x[29..0]"
// Retrieval info: USED_PORT: data47x 0 0 30 0 INPUT NODEFVAL "data47x[29..0]"
// Retrieval info: USED_PORT: data48x 0 0 30 0 INPUT NODEFVAL "data48x[29..0]"
// Retrieval info: USED_PORT: data49x 0 0 30 0 INPUT NODEFVAL "data49x[29..0]"
// Retrieval info: USED_PORT: data4x 0 0 30 0 INPUT NODEFVAL "data4x[29..0]"
// Retrieval info: USED_PORT: data50x 0 0 30 0 INPUT NODEFVAL "data50x[29..0]"
// Retrieval info: USED_PORT: data51x 0 0 30 0 INPUT NODEFVAL "data51x[29..0]"
// Retrieval info: USED_PORT: data52x 0 0 30 0 INPUT NODEFVAL "data52x[29..0]"
// Retrieval info: USED_PORT: data53x 0 0 30 0 INPUT NODEFVAL "data53x[29..0]"
// Retrieval info: USED_PORT: data54x 0 0 30 0 INPUT NODEFVAL "data54x[29..0]"
// Retrieval info: USED_PORT: data55x 0 0 30 0 INPUT NODEFVAL "data55x[29..0]"
// Retrieval info: USED_PORT: data56x 0 0 30 0 INPUT NODEFVAL "data56x[29..0]"
// Retrieval info: USED_PORT: data57x 0 0 30 0 INPUT NODEFVAL "data57x[29..0]"
// Retrieval info: USED_PORT: data58x 0 0 30 0 INPUT NODEFVAL "data58x[29..0]"
// Retrieval info: USED_PORT: data59x 0 0 30 0 INPUT NODEFVAL "data59x[29..0]"
// Retrieval info: USED_PORT: data5x 0 0 30 0 INPUT NODEFVAL "data5x[29..0]"
// Retrieval info: USED_PORT: data60x 0 0 30 0 INPUT NODEFVAL "data60x[29..0]"
// Retrieval info: USED_PORT: data61x 0 0 30 0 INPUT NODEFVAL "data61x[29..0]"
// Retrieval info: USED_PORT: data62x 0 0 30 0 INPUT NODEFVAL "data62x[29..0]"
// Retrieval info: USED_PORT: data63x 0 0 30 0 INPUT NODEFVAL "data63x[29..0]"
// Retrieval info: USED_PORT: data64x 0 0 30 0 INPUT NODEFVAL "data64x[29..0]"
// Retrieval info: USED_PORT: data65x 0 0 30 0 INPUT NODEFVAL "data65x[29..0]"
// Retrieval info: USED_PORT: data66x 0 0 30 0 INPUT NODEFVAL "data66x[29..0]"
// Retrieval info: USED_PORT: data67x 0 0 30 0 INPUT NODEFVAL "data67x[29..0]"
// Retrieval info: USED_PORT: data68x 0 0 30 0 INPUT NODEFVAL "data68x[29..0]"
// Retrieval info: USED_PORT: data69x 0 0 30 0 INPUT NODEFVAL "data69x[29..0]"
// Retrieval info: USED_PORT: data6x 0 0 30 0 INPUT NODEFVAL "data6x[29..0]"
// Retrieval info: USED_PORT: data70x 0 0 30 0 INPUT NODEFVAL "data70x[29..0]"
// Retrieval info: USED_PORT: data71x 0 0 30 0 INPUT NODEFVAL "data71x[29..0]"
// Retrieval info: USED_PORT: data72x 0 0 30 0 INPUT NODEFVAL "data72x[29..0]"
// Retrieval info: USED_PORT: data73x 0 0 30 0 INPUT NODEFVAL "data73x[29..0]"
// Retrieval info: USED_PORT: data74x 0 0 30 0 INPUT NODEFVAL "data74x[29..0]"
// Retrieval info: USED_PORT: data75x 0 0 30 0 INPUT NODEFVAL "data75x[29..0]"
// Retrieval info: USED_PORT: data76x 0 0 30 0 INPUT NODEFVAL "data76x[29..0]"
// Retrieval info: USED_PORT: data77x 0 0 30 0 INPUT NODEFVAL "data77x[29..0]"
// Retrieval info: USED_PORT: data78x 0 0 30 0 INPUT NODEFVAL "data78x[29..0]"
// Retrieval info: USED_PORT: data79x 0 0 30 0 INPUT NODEFVAL "data79x[29..0]"
// Retrieval info: USED_PORT: data7x 0 0 30 0 INPUT NODEFVAL "data7x[29..0]"
// Retrieval info: USED_PORT: data8x 0 0 30 0 INPUT NODEFVAL "data8x[29..0]"
// Retrieval info: USED_PORT: data9x 0 0 30 0 INPUT NODEFVAL "data9x[29..0]"
// Retrieval info: USED_PORT: result 0 0 37 0 OUTPUT NODEFVAL "result[36..0]"
// Retrieval info: CONNECT: @data 0 0 30 0 data0x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 300 data10x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 330 data11x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 360 data12x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 390 data13x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 420 data14x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 450 data15x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 480 data16x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 510 data17x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 540 data18x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 570 data19x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 30 data1x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 600 data20x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 630 data21x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 660 data22x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 690 data23x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 720 data24x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 750 data25x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 780 data26x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 810 data27x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 840 data28x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 870 data29x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 60 data2x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 900 data30x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 930 data31x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 960 data32x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 990 data33x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1020 data34x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1050 data35x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1080 data36x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1110 data37x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1140 data38x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1170 data39x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 90 data3x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1200 data40x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1230 data41x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1260 data42x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1290 data43x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1320 data44x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1350 data45x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1380 data46x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1410 data47x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1440 data48x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1470 data49x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 120 data4x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1500 data50x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1530 data51x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1560 data52x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1590 data53x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1620 data54x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1650 data55x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1680 data56x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1710 data57x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1740 data58x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1770 data59x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 150 data5x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1800 data60x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1830 data61x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1860 data62x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1890 data63x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1920 data64x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1950 data65x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 1980 data66x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 2010 data67x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 2040 data68x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 2070 data69x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 180 data6x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 2100 data70x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 2130 data71x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 2160 data72x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 2190 data73x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 2220 data74x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 2250 data75x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 2280 data76x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 2310 data77x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 2340 data78x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 2370 data79x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 210 data7x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 240 data8x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 270 data9x 0 0 30 0
// Retrieval info: CONNECT: result 0 0 37 0 @result 0 0 37 0
// Retrieval info: GEN_FILE: TYPE_NORMAL pAdd_80.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL pAdd_80.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL pAdd_80.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL pAdd_80.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL pAdd_80_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL pAdd_80_bb.v FALSE
// Retrieval info: LIB_FILE: altera_mf
